module MIPS_Testbench ();
reg CLK;
reg RST;
wire CS;
wire WE;
wire [31:0] Mem_Bus;
wire [31:0] Address;
    initial
    begin
        CLK = 0;
    end
        MIPS CPU(CLK, RST, CS, WE, Address, Mem_Bus);
        Memory MEM(CS, WE, CLK, Address, Mem_Bus);
    always
    begin
        #10 CLK = !CLK;
    end
    always
    begin
        RST <= 1'b1; //reset the processor
        //Notice that the memory is initialize in the in the memory module not here
        @(posedge CLK);
        // driving reset low here puts processor in normal operating mode
        RST = 1'b0;
        /* add your testing code here */
        // you can add in a 'Halt' signal here as well to test Halt operation 
        // you will be verifying your program operation using the 
// waveform viewer and/or self-checking operations
    $display("TEST COMPLETE");
    $stop;
    end
endmodule
